magic
tech sky130A
magscale 1 2
timestamp 1669384289
<< obsli1 >>
rect 1104 2159 133584 134385
<< obsm1 >>
rect 14 1844 134030 134904
<< metal2 >>
rect 662 136108 718 136708
rect 3882 136108 3938 136708
rect 6458 136108 6514 136708
rect 9678 136108 9734 136708
rect 12254 136108 12310 136708
rect 14830 136108 14886 136708
rect 18050 136108 18106 136708
rect 20626 136108 20682 136708
rect 23846 136108 23902 136708
rect 26422 136108 26478 136708
rect 29642 136108 29698 136708
rect 32218 136108 32274 136708
rect 34794 136108 34850 136708
rect 38014 136108 38070 136708
rect 40590 136108 40646 136708
rect 43810 136108 43866 136708
rect 46386 136108 46442 136708
rect 49606 136108 49662 136708
rect 52182 136108 52238 136708
rect 54758 136108 54814 136708
rect 57978 136108 58034 136708
rect 60554 136108 60610 136708
rect 63774 136108 63830 136708
rect 66350 136108 66406 136708
rect 69570 136108 69626 136708
rect 72146 136108 72202 136708
rect 74722 136108 74778 136708
rect 77942 136108 77998 136708
rect 80518 136108 80574 136708
rect 83738 136108 83794 136708
rect 86314 136108 86370 136708
rect 89534 136108 89590 136708
rect 92110 136108 92166 136708
rect 94686 136108 94742 136708
rect 97906 136108 97962 136708
rect 100482 136108 100538 136708
rect 103702 136108 103758 136708
rect 106278 136108 106334 136708
rect 109498 136108 109554 136708
rect 112074 136108 112130 136708
rect 114650 136108 114706 136708
rect 117870 136108 117926 136708
rect 120446 136108 120502 136708
rect 123666 136108 123722 136708
rect 126242 136108 126298 136708
rect 129462 136108 129518 136708
rect 132038 136108 132094 136708
rect 18 200 74 800
rect 2594 200 2650 800
rect 5170 200 5226 800
rect 8390 200 8446 800
rect 10966 200 11022 800
rect 14186 200 14242 800
rect 16762 200 16818 800
rect 19982 200 20038 800
rect 22558 200 22614 800
rect 25134 200 25190 800
rect 28354 200 28410 800
rect 30930 200 30986 800
rect 34150 200 34206 800
rect 36726 200 36782 800
rect 39946 200 40002 800
rect 42522 200 42578 800
rect 45098 200 45154 800
rect 48318 200 48374 800
rect 50894 200 50950 800
rect 54114 200 54170 800
rect 56690 200 56746 800
rect 59910 200 59966 800
rect 62486 200 62542 800
rect 65062 200 65118 800
rect 68282 200 68338 800
rect 70858 200 70914 800
rect 74078 200 74134 800
rect 76654 200 76710 800
rect 79874 200 79930 800
rect 82450 200 82506 800
rect 85026 200 85082 800
rect 88246 200 88302 800
rect 90822 200 90878 800
rect 94042 200 94098 800
rect 96618 200 96674 800
rect 99838 200 99894 800
rect 102414 200 102470 800
rect 104990 200 105046 800
rect 108210 200 108266 800
rect 110786 200 110842 800
rect 114006 200 114062 800
rect 116582 200 116638 800
rect 119802 200 119858 800
rect 122378 200 122434 800
rect 124954 200 125010 800
rect 128174 200 128230 800
rect 130750 200 130806 800
rect 133970 200 134026 800
<< obsm2 >>
rect 20 136764 134024 136785
rect 20 136052 606 136764
rect 774 136052 3826 136764
rect 3994 136052 6402 136764
rect 6570 136052 9622 136764
rect 9790 136052 12198 136764
rect 12366 136052 14774 136764
rect 14942 136052 17994 136764
rect 18162 136052 20570 136764
rect 20738 136052 23790 136764
rect 23958 136052 26366 136764
rect 26534 136052 29586 136764
rect 29754 136052 32162 136764
rect 32330 136052 34738 136764
rect 34906 136052 37958 136764
rect 38126 136052 40534 136764
rect 40702 136052 43754 136764
rect 43922 136052 46330 136764
rect 46498 136052 49550 136764
rect 49718 136052 52126 136764
rect 52294 136052 54702 136764
rect 54870 136052 57922 136764
rect 58090 136052 60498 136764
rect 60666 136052 63718 136764
rect 63886 136052 66294 136764
rect 66462 136052 69514 136764
rect 69682 136052 72090 136764
rect 72258 136052 74666 136764
rect 74834 136052 77886 136764
rect 78054 136052 80462 136764
rect 80630 136052 83682 136764
rect 83850 136052 86258 136764
rect 86426 136052 89478 136764
rect 89646 136052 92054 136764
rect 92222 136052 94630 136764
rect 94798 136052 97850 136764
rect 98018 136052 100426 136764
rect 100594 136052 103646 136764
rect 103814 136052 106222 136764
rect 106390 136052 109442 136764
rect 109610 136052 112018 136764
rect 112186 136052 114594 136764
rect 114762 136052 117814 136764
rect 117982 136052 120390 136764
rect 120558 136052 123610 136764
rect 123778 136052 126186 136764
rect 126354 136052 129406 136764
rect 129574 136052 131982 136764
rect 132150 136052 134024 136764
rect 20 856 134024 136052
rect 130 800 2538 856
rect 2706 800 5114 856
rect 5282 800 8334 856
rect 8502 800 10910 856
rect 11078 800 14130 856
rect 14298 800 16706 856
rect 16874 800 19926 856
rect 20094 800 22502 856
rect 22670 800 25078 856
rect 25246 800 28298 856
rect 28466 800 30874 856
rect 31042 800 34094 856
rect 34262 800 36670 856
rect 36838 800 39890 856
rect 40058 800 42466 856
rect 42634 800 45042 856
rect 45210 800 48262 856
rect 48430 800 50838 856
rect 51006 800 54058 856
rect 54226 800 56634 856
rect 56802 800 59854 856
rect 60022 800 62430 856
rect 62598 800 65006 856
rect 65174 800 68226 856
rect 68394 800 70802 856
rect 70970 800 74022 856
rect 74190 800 76598 856
rect 76766 800 79818 856
rect 79986 800 82394 856
rect 82562 800 84970 856
rect 85138 800 88190 856
rect 88358 800 90766 856
rect 90934 800 93986 856
rect 94154 800 96562 856
rect 96730 800 99782 856
rect 99950 800 102358 856
rect 102526 800 104934 856
rect 105102 800 108154 856
rect 108322 800 110730 856
rect 110898 800 113950 856
rect 114118 800 116526 856
rect 116694 800 119746 856
rect 119914 800 122322 856
rect 122490 800 124898 856
rect 125066 800 128118 856
rect 128286 800 130694 856
rect 130862 800 133914 856
<< metal3 >>
rect 133964 136688 134564 136808
rect 200 135328 800 135448
rect 133964 133968 134564 134088
rect 200 131928 800 132048
rect 133964 131248 134564 131368
rect 200 129208 800 129328
rect 133964 127848 134564 127968
rect 200 126488 800 126608
rect 133964 125128 134564 125248
rect 200 123088 800 123208
rect 133964 121728 134564 121848
rect 200 120368 800 120488
rect 133964 119008 134564 119128
rect 200 116968 800 117088
rect 133964 115608 134564 115728
rect 200 114248 800 114368
rect 133964 112888 134564 113008
rect 200 110848 800 110968
rect 133964 110168 134564 110288
rect 200 108128 800 108248
rect 133964 106768 134564 106888
rect 200 105408 800 105528
rect 133964 104048 134564 104168
rect 200 102008 800 102128
rect 133964 100648 134564 100768
rect 200 99288 800 99408
rect 133964 97928 134564 98048
rect 200 95888 800 96008
rect 133964 94528 134564 94648
rect 200 93168 800 93288
rect 133964 91808 134564 91928
rect 200 89768 800 89888
rect 133964 89088 134564 89208
rect 200 87048 800 87168
rect 133964 85688 134564 85808
rect 200 84328 800 84448
rect 133964 82968 134564 83088
rect 200 80928 800 81048
rect 133964 79568 134564 79688
rect 200 78208 800 78328
rect 133964 76848 134564 76968
rect 200 74808 800 74928
rect 133964 73448 134564 73568
rect 200 72088 800 72208
rect 133964 70728 134564 70848
rect 200 68688 800 68808
rect 133964 68008 134564 68128
rect 200 65968 800 66088
rect 133964 64608 134564 64728
rect 200 63248 800 63368
rect 133964 61888 134564 62008
rect 200 59848 800 59968
rect 133964 58488 134564 58608
rect 200 57128 800 57248
rect 133964 55768 134564 55888
rect 200 53728 800 53848
rect 133964 52368 134564 52488
rect 200 51008 800 51128
rect 133964 49648 134564 49768
rect 200 47608 800 47728
rect 133964 46928 134564 47048
rect 200 44888 800 45008
rect 133964 43528 134564 43648
rect 200 42168 800 42288
rect 133964 40808 134564 40928
rect 200 38768 800 38888
rect 133964 37408 134564 37528
rect 200 36048 800 36168
rect 133964 34688 134564 34808
rect 200 32648 800 32768
rect 133964 31288 134564 31408
rect 200 29928 800 30048
rect 133964 28568 134564 28688
rect 200 26528 800 26648
rect 133964 25848 134564 25968
rect 200 23808 800 23928
rect 133964 22448 134564 22568
rect 200 21088 800 21208
rect 133964 19728 134564 19848
rect 200 17688 800 17808
rect 133964 16328 134564 16448
rect 200 14968 800 15088
rect 133964 13608 134564 13728
rect 200 11568 800 11688
rect 133964 10208 134564 10328
rect 200 8848 800 8968
rect 133964 7488 134564 7608
rect 200 5448 800 5568
rect 133964 4768 134564 4888
rect 200 2728 800 2848
rect 133964 1368 134564 1488
<< obsm3 >>
rect 800 136608 133884 136781
rect 800 135528 133964 136608
rect 880 135248 133964 135528
rect 800 134168 133964 135248
rect 800 133888 133884 134168
rect 800 132128 133964 133888
rect 880 131848 133964 132128
rect 800 131448 133964 131848
rect 800 131168 133884 131448
rect 800 129408 133964 131168
rect 880 129128 133964 129408
rect 800 128048 133964 129128
rect 800 127768 133884 128048
rect 800 126688 133964 127768
rect 880 126408 133964 126688
rect 800 125328 133964 126408
rect 800 125048 133884 125328
rect 800 123288 133964 125048
rect 880 123008 133964 123288
rect 800 121928 133964 123008
rect 800 121648 133884 121928
rect 800 120568 133964 121648
rect 880 120288 133964 120568
rect 800 119208 133964 120288
rect 800 118928 133884 119208
rect 800 117168 133964 118928
rect 880 116888 133964 117168
rect 800 115808 133964 116888
rect 800 115528 133884 115808
rect 800 114448 133964 115528
rect 880 114168 133964 114448
rect 800 113088 133964 114168
rect 800 112808 133884 113088
rect 800 111048 133964 112808
rect 880 110768 133964 111048
rect 800 110368 133964 110768
rect 800 110088 133884 110368
rect 800 108328 133964 110088
rect 880 108048 133964 108328
rect 800 106968 133964 108048
rect 800 106688 133884 106968
rect 800 105608 133964 106688
rect 880 105328 133964 105608
rect 800 104248 133964 105328
rect 800 103968 133884 104248
rect 800 102208 133964 103968
rect 880 101928 133964 102208
rect 800 100848 133964 101928
rect 800 100568 133884 100848
rect 800 99488 133964 100568
rect 880 99208 133964 99488
rect 800 98128 133964 99208
rect 800 97848 133884 98128
rect 800 96088 133964 97848
rect 880 95808 133964 96088
rect 800 94728 133964 95808
rect 800 94448 133884 94728
rect 800 93368 133964 94448
rect 880 93088 133964 93368
rect 800 92008 133964 93088
rect 800 91728 133884 92008
rect 800 89968 133964 91728
rect 880 89688 133964 89968
rect 800 89288 133964 89688
rect 800 89008 133884 89288
rect 800 87248 133964 89008
rect 880 86968 133964 87248
rect 800 85888 133964 86968
rect 800 85608 133884 85888
rect 800 84528 133964 85608
rect 880 84248 133964 84528
rect 800 83168 133964 84248
rect 800 82888 133884 83168
rect 800 81128 133964 82888
rect 880 80848 133964 81128
rect 800 79768 133964 80848
rect 800 79488 133884 79768
rect 800 78408 133964 79488
rect 880 78128 133964 78408
rect 800 77048 133964 78128
rect 800 76768 133884 77048
rect 800 75008 133964 76768
rect 880 74728 133964 75008
rect 800 73648 133964 74728
rect 800 73368 133884 73648
rect 800 72288 133964 73368
rect 880 72008 133964 72288
rect 800 70928 133964 72008
rect 800 70648 133884 70928
rect 800 68888 133964 70648
rect 880 68608 133964 68888
rect 800 68208 133964 68608
rect 800 67928 133884 68208
rect 800 66168 133964 67928
rect 880 65888 133964 66168
rect 800 64808 133964 65888
rect 800 64528 133884 64808
rect 800 63448 133964 64528
rect 880 63168 133964 63448
rect 800 62088 133964 63168
rect 800 61808 133884 62088
rect 800 60048 133964 61808
rect 880 59768 133964 60048
rect 800 58688 133964 59768
rect 800 58408 133884 58688
rect 800 57328 133964 58408
rect 880 57048 133964 57328
rect 800 55968 133964 57048
rect 800 55688 133884 55968
rect 800 53928 133964 55688
rect 880 53648 133964 53928
rect 800 52568 133964 53648
rect 800 52288 133884 52568
rect 800 51208 133964 52288
rect 880 50928 133964 51208
rect 800 49848 133964 50928
rect 800 49568 133884 49848
rect 800 47808 133964 49568
rect 880 47528 133964 47808
rect 800 47128 133964 47528
rect 800 46848 133884 47128
rect 800 45088 133964 46848
rect 880 44808 133964 45088
rect 800 43728 133964 44808
rect 800 43448 133884 43728
rect 800 42368 133964 43448
rect 880 42088 133964 42368
rect 800 41008 133964 42088
rect 800 40728 133884 41008
rect 800 38968 133964 40728
rect 880 38688 133964 38968
rect 800 37608 133964 38688
rect 800 37328 133884 37608
rect 800 36248 133964 37328
rect 880 35968 133964 36248
rect 800 34888 133964 35968
rect 800 34608 133884 34888
rect 800 32848 133964 34608
rect 880 32568 133964 32848
rect 800 31488 133964 32568
rect 800 31208 133884 31488
rect 800 30128 133964 31208
rect 880 29848 133964 30128
rect 800 28768 133964 29848
rect 800 28488 133884 28768
rect 800 26728 133964 28488
rect 880 26448 133964 26728
rect 800 26048 133964 26448
rect 800 25768 133884 26048
rect 800 24008 133964 25768
rect 880 23728 133964 24008
rect 800 22648 133964 23728
rect 800 22368 133884 22648
rect 800 21288 133964 22368
rect 880 21008 133964 21288
rect 800 19928 133964 21008
rect 800 19648 133884 19928
rect 800 17888 133964 19648
rect 880 17608 133964 17888
rect 800 16528 133964 17608
rect 800 16248 133884 16528
rect 800 15168 133964 16248
rect 880 14888 133964 15168
rect 800 13808 133964 14888
rect 800 13528 133884 13808
rect 800 11768 133964 13528
rect 880 11488 133964 11768
rect 800 10408 133964 11488
rect 800 10128 133884 10408
rect 800 9048 133964 10128
rect 880 8768 133964 9048
rect 800 7688 133964 8768
rect 800 7408 133884 7688
rect 800 5648 133964 7408
rect 880 5368 133964 5648
rect 800 4968 133964 5368
rect 800 4688 133884 4968
rect 800 2928 133964 4688
rect 880 2648 133964 2928
rect 800 1568 133964 2648
rect 800 1395 133884 1568
<< metal4 >>
rect 4208 2128 4528 134416
rect 19568 2128 19888 134416
rect 34928 2128 35248 134416
rect 50288 2128 50608 134416
rect 65648 2128 65968 134416
rect 81008 2128 81328 134416
rect 96368 2128 96688 134416
rect 111728 2128 112048 134416
rect 127088 2128 127408 134416
<< obsm4 >>
rect 8155 2048 19488 134197
rect 19968 2048 34848 134197
rect 35328 2048 50208 134197
rect 50688 2048 65568 134197
rect 66048 2048 80928 134197
rect 81408 2048 96288 134197
rect 96768 2048 111648 134197
rect 112128 2048 122669 134197
rect 8155 1803 122669 2048
<< labels >>
rlabel metal2 s 65062 200 65118 800 6 dbg_freeze_i
port 1 nsew signal input
rlabel metal3 s 133964 133968 134564 134088 6 irq_gfx_o
port 2 nsew signal output
rlabel metal3 s 200 126488 800 126608 6 lt24_cs_n_o
port 3 nsew signal output
rlabel metal3 s 200 29928 800 30048 6 lt24_d_en_o
port 4 nsew signal output
rlabel metal2 s 10966 200 11022 800 6 lt24_d_i[0]
port 5 nsew signal input
rlabel metal2 s 114006 200 114062 800 6 lt24_d_i[10]
port 6 nsew signal input
rlabel metal3 s 200 129208 800 129328 6 lt24_d_i[11]
port 7 nsew signal input
rlabel metal2 s 36726 200 36782 800 6 lt24_d_i[12]
port 8 nsew signal input
rlabel metal3 s 133964 13608 134564 13728 6 lt24_d_i[13]
port 9 nsew signal input
rlabel metal3 s 200 5448 800 5568 6 lt24_d_i[14]
port 10 nsew signal input
rlabel metal3 s 133964 31288 134564 31408 6 lt24_d_i[15]
port 11 nsew signal input
rlabel metal2 s 119802 200 119858 800 6 lt24_d_i[1]
port 12 nsew signal input
rlabel metal2 s 43810 136108 43866 136708 6 lt24_d_i[2]
port 13 nsew signal input
rlabel metal3 s 200 51008 800 51128 6 lt24_d_i[3]
port 14 nsew signal input
rlabel metal3 s 200 65968 800 66088 6 lt24_d_i[4]
port 15 nsew signal input
rlabel metal2 s 74722 136108 74778 136708 6 lt24_d_i[5]
port 16 nsew signal input
rlabel metal2 s 30930 200 30986 800 6 lt24_d_i[6]
port 17 nsew signal input
rlabel metal2 s 38014 136108 38070 136708 6 lt24_d_i[7]
port 18 nsew signal input
rlabel metal3 s 200 68688 800 68808 6 lt24_d_i[8]
port 19 nsew signal input
rlabel metal3 s 200 57128 800 57248 6 lt24_d_i[9]
port 20 nsew signal input
rlabel metal2 s 88246 200 88302 800 6 lt24_d_o[0]
port 21 nsew signal output
rlabel metal2 s 120446 136108 120502 136708 6 lt24_d_o[10]
port 22 nsew signal output
rlabel metal2 s 72146 136108 72202 136708 6 lt24_d_o[11]
port 23 nsew signal output
rlabel metal3 s 200 78208 800 78328 6 lt24_d_o[12]
port 24 nsew signal output
rlabel metal3 s 133964 34688 134564 34808 6 lt24_d_o[13]
port 25 nsew signal output
rlabel metal2 s 26422 136108 26478 136708 6 lt24_d_o[14]
port 26 nsew signal output
rlabel metal3 s 133964 79568 134564 79688 6 lt24_d_o[15]
port 27 nsew signal output
rlabel metal3 s 200 123088 800 123208 6 lt24_d_o[1]
port 28 nsew signal output
rlabel metal2 s 117870 136108 117926 136708 6 lt24_d_o[2]
port 29 nsew signal output
rlabel metal2 s 83738 136108 83794 136708 6 lt24_d_o[3]
port 30 nsew signal output
rlabel metal3 s 200 89768 800 89888 6 lt24_d_o[4]
port 31 nsew signal output
rlabel metal3 s 133964 115608 134564 115728 6 lt24_d_o[5]
port 32 nsew signal output
rlabel metal3 s 133964 100648 134564 100768 6 lt24_d_o[6]
port 33 nsew signal output
rlabel metal2 s 128174 200 128230 800 6 lt24_d_o[7]
port 34 nsew signal output
rlabel metal3 s 200 32648 800 32768 6 lt24_d_o[8]
port 35 nsew signal output
rlabel metal2 s 40590 136108 40646 136708 6 lt24_d_o[9]
port 36 nsew signal output
rlabel metal3 s 133964 104048 134564 104168 6 lt24_on_o
port 37 nsew signal output
rlabel metal3 s 200 59848 800 59968 6 lt24_rd_n_o
port 38 nsew signal output
rlabel metal3 s 133964 16328 134564 16448 6 lt24_reset_n_o
port 39 nsew signal output
rlabel metal3 s 133964 97928 134564 98048 6 lt24_rs_o
port 40 nsew signal output
rlabel metal3 s 133964 40808 134564 40928 6 lt24_wr_n_o
port 41 nsew signal output
rlabel metal2 s 103702 136108 103758 136708 6 lut_ram_addr_o[0]
port 42 nsew signal output
rlabel metal2 s 100482 136108 100538 136708 6 lut_ram_addr_o[1]
port 43 nsew signal output
rlabel metal3 s 133964 121728 134564 121848 6 lut_ram_addr_o[2]
port 44 nsew signal output
rlabel metal3 s 200 95888 800 96008 6 lut_ram_addr_o[3]
port 45 nsew signal output
rlabel metal2 s 29642 136108 29698 136708 6 lut_ram_addr_o[4]
port 46 nsew signal output
rlabel metal2 s 54114 200 54170 800 6 lut_ram_addr_o[5]
port 47 nsew signal output
rlabel metal3 s 133964 131248 134564 131368 6 lut_ram_addr_o[6]
port 48 nsew signal output
rlabel metal3 s 200 84328 800 84448 6 lut_ram_addr_o[7]
port 49 nsew signal output
rlabel metal3 s 200 2728 800 2848 6 lut_ram_addr_o[8]
port 50 nsew signal output
rlabel metal2 s 22558 200 22614 800 6 lut_ram_cen_o
port 51 nsew signal output
rlabel metal3 s 133964 73448 134564 73568 6 lut_ram_din_o[0]
port 52 nsew signal output
rlabel metal3 s 133964 19728 134564 19848 6 lut_ram_din_o[10]
port 53 nsew signal output
rlabel metal2 s 54758 136108 54814 136708 6 lut_ram_din_o[11]
port 54 nsew signal output
rlabel metal2 s 42522 200 42578 800 6 lut_ram_din_o[12]
port 55 nsew signal output
rlabel metal2 s 85026 200 85082 800 6 lut_ram_din_o[13]
port 56 nsew signal output
rlabel metal2 s 662 136108 718 136708 6 lut_ram_din_o[14]
port 57 nsew signal output
rlabel metal3 s 133964 119008 134564 119128 6 lut_ram_din_o[15]
port 58 nsew signal output
rlabel metal3 s 133964 61888 134564 62008 6 lut_ram_din_o[1]
port 59 nsew signal output
rlabel metal2 s 49606 136108 49662 136708 6 lut_ram_din_o[2]
port 60 nsew signal output
rlabel metal2 s 99838 200 99894 800 6 lut_ram_din_o[3]
port 61 nsew signal output
rlabel metal2 s 106278 136108 106334 136708 6 lut_ram_din_o[4]
port 62 nsew signal output
rlabel metal3 s 200 72088 800 72208 6 lut_ram_din_o[5]
port 63 nsew signal output
rlabel metal2 s 126242 136108 126298 136708 6 lut_ram_din_o[6]
port 64 nsew signal output
rlabel metal3 s 133964 1368 134564 1488 6 lut_ram_din_o[7]
port 65 nsew signal output
rlabel metal2 s 123666 136108 123722 136708 6 lut_ram_din_o[8]
port 66 nsew signal output
rlabel metal3 s 133964 25848 134564 25968 6 lut_ram_din_o[9]
port 67 nsew signal output
rlabel metal2 s 62486 200 62542 800 6 lut_ram_dout_i[0]
port 68 nsew signal input
rlabel metal3 s 133964 55768 134564 55888 6 lut_ram_dout_i[10]
port 69 nsew signal input
rlabel metal2 s 112074 136108 112130 136708 6 lut_ram_dout_i[11]
port 70 nsew signal input
rlabel metal2 s 102414 200 102470 800 6 lut_ram_dout_i[12]
port 71 nsew signal input
rlabel metal2 s 39946 200 40002 800 6 lut_ram_dout_i[13]
port 72 nsew signal input
rlabel metal3 s 200 17688 800 17808 6 lut_ram_dout_i[14]
port 73 nsew signal input
rlabel metal3 s 200 131928 800 132048 6 lut_ram_dout_i[15]
port 74 nsew signal input
rlabel metal3 s 200 53728 800 53848 6 lut_ram_dout_i[1]
port 75 nsew signal input
rlabel metal3 s 133964 68008 134564 68128 6 lut_ram_dout_i[2]
port 76 nsew signal input
rlabel metal2 s 52182 136108 52238 136708 6 lut_ram_dout_i[3]
port 77 nsew signal input
rlabel metal3 s 200 99288 800 99408 6 lut_ram_dout_i[4]
port 78 nsew signal input
rlabel metal2 s 14830 136108 14886 136708 6 lut_ram_dout_i[5]
port 79 nsew signal input
rlabel metal3 s 133964 110168 134564 110288 6 lut_ram_dout_i[6]
port 80 nsew signal input
rlabel metal2 s 6458 136108 6514 136708 6 lut_ram_dout_i[7]
port 81 nsew signal input
rlabel metal2 s 32218 136108 32274 136708 6 lut_ram_dout_i[8]
port 82 nsew signal input
rlabel metal2 s 104990 200 105046 800 6 lut_ram_dout_i[9]
port 83 nsew signal input
rlabel metal2 s 69570 136108 69626 136708 6 lut_ram_wen_o
port 84 nsew signal output
rlabel metal2 s 132038 136108 132094 136708 6 mclk
port 85 nsew signal input
rlabel metal3 s 200 74808 800 74928 6 per_addr_i[0]
port 86 nsew signal input
rlabel metal2 s 5170 200 5226 800 6 per_addr_i[10]
port 87 nsew signal input
rlabel metal2 s 45098 200 45154 800 6 per_addr_i[11]
port 88 nsew signal input
rlabel metal2 s 23846 136108 23902 136708 6 per_addr_i[12]
port 89 nsew signal input
rlabel metal3 s 133964 4768 134564 4888 6 per_addr_i[13]
port 90 nsew signal input
rlabel metal2 s 50894 200 50950 800 6 per_addr_i[1]
port 91 nsew signal input
rlabel metal3 s 200 21088 800 21208 6 per_addr_i[2]
port 92 nsew signal input
rlabel metal2 s 110786 200 110842 800 6 per_addr_i[3]
port 93 nsew signal input
rlabel metal2 s 82450 200 82506 800 6 per_addr_i[4]
port 94 nsew signal input
rlabel metal3 s 133964 70728 134564 70848 6 per_addr_i[5]
port 95 nsew signal input
rlabel metal3 s 133964 46928 134564 47048 6 per_addr_i[6]
port 96 nsew signal input
rlabel metal2 s 114650 136108 114706 136708 6 per_addr_i[7]
port 97 nsew signal input
rlabel metal2 s 86314 136108 86370 136708 6 per_addr_i[8]
port 98 nsew signal input
rlabel metal2 s 108210 200 108266 800 6 per_addr_i[9]
port 99 nsew signal input
rlabel metal3 s 133964 127848 134564 127968 6 per_din_i[0]
port 100 nsew signal input
rlabel metal3 s 200 8848 800 8968 6 per_din_i[10]
port 101 nsew signal input
rlabel metal3 s 200 44888 800 45008 6 per_din_i[11]
port 102 nsew signal input
rlabel metal2 s 46386 136108 46442 136708 6 per_din_i[12]
port 103 nsew signal input
rlabel metal2 s 3882 136108 3938 136708 6 per_din_i[13]
port 104 nsew signal input
rlabel metal3 s 200 110848 800 110968 6 per_din_i[14]
port 105 nsew signal input
rlabel metal2 s 12254 136108 12310 136708 6 per_din_i[15]
port 106 nsew signal input
rlabel metal3 s 133964 76848 134564 76968 6 per_din_i[1]
port 107 nsew signal input
rlabel metal2 s 133970 200 134026 800 6 per_din_i[2]
port 108 nsew signal input
rlabel metal3 s 200 14968 800 15088 6 per_din_i[3]
port 109 nsew signal input
rlabel metal3 s 133964 82968 134564 83088 6 per_din_i[4]
port 110 nsew signal input
rlabel metal2 s 70858 200 70914 800 6 per_din_i[5]
port 111 nsew signal input
rlabel metal3 s 200 38768 800 38888 6 per_din_i[6]
port 112 nsew signal input
rlabel metal2 s 57978 136108 58034 136708 6 per_din_i[7]
port 113 nsew signal input
rlabel metal2 s 96618 200 96674 800 6 per_din_i[8]
port 114 nsew signal input
rlabel metal2 s 124954 200 125010 800 6 per_din_i[9]
port 115 nsew signal input
rlabel metal3 s 200 102008 800 102128 6 per_dout_o[0]
port 116 nsew signal output
rlabel metal3 s 133964 52368 134564 52488 6 per_dout_o[10]
port 117 nsew signal output
rlabel metal2 s 60554 136108 60610 136708 6 per_dout_o[11]
port 118 nsew signal output
rlabel metal2 s 80518 136108 80574 136708 6 per_dout_o[12]
port 119 nsew signal output
rlabel metal2 s 77942 136108 77998 136708 6 per_dout_o[13]
port 120 nsew signal output
rlabel metal3 s 200 108128 800 108248 6 per_dout_o[14]
port 121 nsew signal output
rlabel metal2 s 19982 200 20038 800 6 per_dout_o[15]
port 122 nsew signal output
rlabel metal3 s 133964 22448 134564 22568 6 per_dout_o[1]
port 123 nsew signal output
rlabel metal2 s 59910 200 59966 800 6 per_dout_o[2]
port 124 nsew signal output
rlabel metal3 s 133964 112888 134564 113008 6 per_dout_o[3]
port 125 nsew signal output
rlabel metal3 s 133964 85688 134564 85808 6 per_dout_o[4]
port 126 nsew signal output
rlabel metal2 s 89534 136108 89590 136708 6 per_dout_o[5]
port 127 nsew signal output
rlabel metal2 s 14186 200 14242 800 6 per_dout_o[6]
port 128 nsew signal output
rlabel metal3 s 133964 37408 134564 37528 6 per_dout_o[7]
port 129 nsew signal output
rlabel metal3 s 200 120368 800 120488 6 per_dout_o[8]
port 130 nsew signal output
rlabel metal2 s 34794 136108 34850 136708 6 per_dout_o[9]
port 131 nsew signal output
rlabel metal3 s 133964 58488 134564 58608 6 per_en_i
port 132 nsew signal input
rlabel metal3 s 133964 7488 134564 7608 6 per_we_i[0]
port 133 nsew signal input
rlabel metal2 s 74078 200 74134 800 6 per_we_i[1]
port 134 nsew signal input
rlabel metal3 s 133964 106768 134564 106888 6 puc_rst
port 135 nsew signal input
rlabel metal4 s 4208 2128 4528 134416 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 134416 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 134416 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 134416 6 vccd1
port 136 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 134416 6 vccd1
port 136 nsew power bidirectional
rlabel metal3 s 200 23808 800 23928 6 vid_ram_addr_o[0]
port 137 nsew signal output
rlabel metal2 s 34150 200 34206 800 6 vid_ram_addr_o[10]
port 138 nsew signal output
rlabel metal3 s 133964 43528 134564 43648 6 vid_ram_addr_o[11]
port 139 nsew signal output
rlabel metal2 s 90822 200 90878 800 6 vid_ram_addr_o[12]
port 140 nsew signal output
rlabel metal3 s 133964 10208 134564 10328 6 vid_ram_addr_o[13]
port 141 nsew signal output
rlabel metal2 s 9678 136108 9734 136708 6 vid_ram_addr_o[14]
port 142 nsew signal output
rlabel metal2 s 116582 200 116638 800 6 vid_ram_addr_o[15]
port 143 nsew signal output
rlabel metal2 s 16762 200 16818 800 6 vid_ram_addr_o[16]
port 144 nsew signal output
rlabel metal2 s 56690 200 56746 800 6 vid_ram_addr_o[1]
port 145 nsew signal output
rlabel metal3 s 200 47608 800 47728 6 vid_ram_addr_o[2]
port 146 nsew signal output
rlabel metal3 s 133964 125128 134564 125248 6 vid_ram_addr_o[3]
port 147 nsew signal output
rlabel metal3 s 133964 89088 134564 89208 6 vid_ram_addr_o[4]
port 148 nsew signal output
rlabel metal2 s 122378 200 122434 800 6 vid_ram_addr_o[5]
port 149 nsew signal output
rlabel metal3 s 200 63248 800 63368 6 vid_ram_addr_o[6]
port 150 nsew signal output
rlabel metal3 s 133964 49648 134564 49768 6 vid_ram_addr_o[7]
port 151 nsew signal output
rlabel metal2 s 2594 200 2650 800 6 vid_ram_addr_o[8]
port 152 nsew signal output
rlabel metal3 s 200 42168 800 42288 6 vid_ram_addr_o[9]
port 153 nsew signal output
rlabel metal3 s 133964 136688 134564 136808 6 vid_ram_cen_o
port 154 nsew signal output
rlabel metal2 s 130750 200 130806 800 6 vid_ram_din_o[0]
port 155 nsew signal output
rlabel metal2 s 129462 136108 129518 136708 6 vid_ram_din_o[10]
port 156 nsew signal output
rlabel metal3 s 200 87048 800 87168 6 vid_ram_din_o[11]
port 157 nsew signal output
rlabel metal3 s 200 93168 800 93288 6 vid_ram_din_o[12]
port 158 nsew signal output
rlabel metal2 s 79874 200 79930 800 6 vid_ram_din_o[13]
port 159 nsew signal output
rlabel metal2 s 18 200 74 800 6 vid_ram_din_o[14]
port 160 nsew signal output
rlabel metal3 s 200 11568 800 11688 6 vid_ram_din_o[15]
port 161 nsew signal output
rlabel metal3 s 200 105408 800 105528 6 vid_ram_din_o[1]
port 162 nsew signal output
rlabel metal2 s 18050 136108 18106 136708 6 vid_ram_din_o[2]
port 163 nsew signal output
rlabel metal2 s 66350 136108 66406 136708 6 vid_ram_din_o[3]
port 164 nsew signal output
rlabel metal3 s 200 80928 800 81048 6 vid_ram_din_o[4]
port 165 nsew signal output
rlabel metal2 s 25134 200 25190 800 6 vid_ram_din_o[5]
port 166 nsew signal output
rlabel metal2 s 8390 200 8446 800 6 vid_ram_din_o[6]
port 167 nsew signal output
rlabel metal2 s 92110 136108 92166 136708 6 vid_ram_din_o[7]
port 168 nsew signal output
rlabel metal2 s 63774 136108 63830 136708 6 vid_ram_din_o[8]
port 169 nsew signal output
rlabel metal2 s 68282 200 68338 800 6 vid_ram_din_o[9]
port 170 nsew signal output
rlabel metal2 s 109498 136108 109554 136708 6 vid_ram_dout_i[0]
port 171 nsew signal input
rlabel metal3 s 133964 28568 134564 28688 6 vid_ram_dout_i[10]
port 172 nsew signal input
rlabel metal3 s 200 114248 800 114368 6 vid_ram_dout_i[11]
port 173 nsew signal input
rlabel metal3 s 133964 94528 134564 94648 6 vid_ram_dout_i[12]
port 174 nsew signal input
rlabel metal2 s 28354 200 28410 800 6 vid_ram_dout_i[13]
port 175 nsew signal input
rlabel metal2 s 48318 200 48374 800 6 vid_ram_dout_i[14]
port 176 nsew signal input
rlabel metal3 s 200 26528 800 26648 6 vid_ram_dout_i[15]
port 177 nsew signal input
rlabel metal3 s 133964 91808 134564 91928 6 vid_ram_dout_i[1]
port 178 nsew signal input
rlabel metal2 s 76654 200 76710 800 6 vid_ram_dout_i[2]
port 179 nsew signal input
rlabel metal2 s 97906 136108 97962 136708 6 vid_ram_dout_i[3]
port 180 nsew signal input
rlabel metal2 s 94686 136108 94742 136708 6 vid_ram_dout_i[4]
port 181 nsew signal input
rlabel metal3 s 200 135328 800 135448 6 vid_ram_dout_i[5]
port 182 nsew signal input
rlabel metal2 s 20626 136108 20682 136708 6 vid_ram_dout_i[6]
port 183 nsew signal input
rlabel metal2 s 94042 200 94098 800 6 vid_ram_dout_i[7]
port 184 nsew signal input
rlabel metal3 s 200 36048 800 36168 6 vid_ram_dout_i[8]
port 185 nsew signal input
rlabel metal3 s 200 116968 800 117088 6 vid_ram_dout_i[9]
port 186 nsew signal input
rlabel metal3 s 133964 64608 134564 64728 6 vid_ram_wen_o
port 187 nsew signal output
rlabel metal4 s 19568 2128 19888 134416 6 vssd1
port 188 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 134416 6 vssd1
port 188 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 134416 6 vssd1
port 188 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 134416 6 vssd1
port 188 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 134764 136908
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 53373872
string GDS_FILE /home/vijayan/CARAVEL_FLOW/mpw7_resubmission/graphics_controller_mpw7/graphics_controller_resubmit/openlane/openGFX430/runs/22_11_25_13_23/results/signoff/openGFX430.magic.gds
string GDS_START 1956040
<< end >>

